module edeco ( 
	e,
	display
	) ;

input [3:0] e;
inout [6:0] display;
