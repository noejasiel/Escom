module multi ( 
	sel,
	a,
	b,
	salida
	) ;

input [1:0] sel;
input [1:0] a;
input [1:0] b;
input [6:0] salida;
