module ff_kjt ( 
	k,
	j,
	t,
	clk,
	q1,
	q2
	) ;

input  k;
input  j;
input  t;
input  clk;
inout  q1;
inout  q2;
