module suma ( 
	c0,
	a1,
	a2,
	a3,
	a4,
	b1,
	b2,
	b3,
	b4,
	s1,
	s2,
	s3,
	s4,
	c1,
	c2,
	c3
	) ;

input  c0;
input  a1;
input  a2;
input  a3;
input  a4;
input  b1;
input  b2;
input  b3;
input  b4;
inout  s1;
inout  s2;
inout  s3;
inout  s4;
inout  c1;
inout  c2;
inout  c3;
