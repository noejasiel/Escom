module sum ( 
	sump,
	sumg,
	salida
	) ;

input [3:0] sump;
input [3:0] sumg;
inout [4:0] salida;
