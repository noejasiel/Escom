module compuertas ( 
	sel,
	a,
	b,
	c,
	salida
	) ;

input [2:0] sel;
input  a;
input  b;
input  c;
inout  salida;
