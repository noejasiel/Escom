module comparadoor ( 
	a,
	b,
	display
	) ;

input [3:0] a;
input [3:0] b;
inout [6:0] display;
