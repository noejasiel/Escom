module ff_rsd ( 
	r,
	s,
	d,
	clk,
	q1,
	q2
	) ;

input  r;
input  s;
input  d;
input  clk;
inout  q1;
inout  q2;
