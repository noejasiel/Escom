module res ( 
	x,
	y,
	s,
	a
	) ;

input  x;
input  y;
inout  s;
inout  a;
