module ff_rsd ( 
	r,
	s,
	d,
	q1,
	q2
	) ;

input  r;
input  s;
input  d;
inout  q1;
inout  q2;
