module and2 ( 
	y0,
	a,
	b,
	c,
	d
	) ;

inout  y0;
input  a;
input  b;
input  c;
input  d;
