module arq_multi ( 
	a,
	b,
	s
	) ;

input [1:0] a;
input [1:0] b;
inout [3:0] s;
