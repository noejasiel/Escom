module suma ( 
	x,
	y,
	z,
	s,
	a
	) ;

input  x;
input  y;
input  z;
inout  s;
inout  a;
