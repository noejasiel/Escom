module multi ( 
	sel,
	b,
	a,
	salida
	) ;

input [1:0] sel;
input [1:0] b;
input [2:0] a;
inout [6:0] salida;
